-- Elementos de Sistemas
-- by Luciano Soares
-- Ram512.vhd

Library ieee;
use ieee.std_logic_1164.all;

entity Ram512 is
	port(
		clock:   in  STD_LOGIC;
		input:   in  STD_LOGIC_VECTOR(15 downto 0);
		load:    in  STD_LOGIC;
		address: in  STD_LOGIC_VECTOR( 8 downto 0);
		output:  out STD_LOGIC_VECTOR(15 downto 0)
	);
end entity;

architecture arch of Ram512 is

	component Ram64 is
		port(
			clock:   in  STD_LOGIC;
			input:   in  STD_LOGIC_VECTOR(15 downto 0);
			load:    in  STD_LOGIC;
			address: in  STD_LOGIC_VECTOR( 5 downto 0);
			output:  out STD_LOGIC_VECTOR(15 downto 0)
		);
	end component;

	component Mux8Way16 is
		port (
				a:   in  STD_LOGIC_VECTOR(15 downto 0);
				b:   in  STD_LOGIC_VECTOR(15 downto 0);
				c:   in  STD_LOGIC_VECTOR(15 downto 0);
				d:   in  STD_LOGIC_VECTOR(15 downto 0);
				e:   in  STD_LOGIC_VECTOR(15 downto 0);
				f:   in  STD_LOGIC_VECTOR(15 downto 0);
				g:   in  STD_LOGIC_VECTOR(15 downto 0);
				h:   in  STD_LOGIC_VECTOR(15 downto 0);
				sel: in  STD_LOGIC_VECTOR( 2 downto 0);
				q:   out STD_LOGIC_VECTOR(15 downto 0));
	end component;

	component DMux8Way is
		port (
			a:   in  STD_LOGIC;
			sel: in  STD_LOGIC_VECTOR(2 downto 0);
			q0:  out STD_LOGIC;
			q1:  out STD_LOGIC;
			q2:  out STD_LOGIC;
			q3:  out STD_LOGIC;
			q4:  out STD_LOGIC;
			q5:  out STD_LOGIC;
			q6:  out STD_LOGIC;
			q7:  out STD_LOGIC);
	end component;

	signal load0, load1, load2, load3, load4, load5, load6, load7 : STD_LOGIC;
	signal output0, output1, output2, output3, output4, output5, output6, output7 : STD_LOGIC_VECTOR(15 downto 0);

begin

	ram0 : Ram64
	port map(
		clock => clock,
		input => input,
		load => load,
		address => address( 5 downto 0),
		output => output
	);
	ram1 : Ram64
	port map(
		clock => clock,
		input => input,
		load => load,
		address => address( 5 downto 0),
		output => output
	);
	ram2 : Ram64
	port map(
		clock => clock,
		input => input,
		load => load,
		address => address( 5 downto 0),
		output => output
	);
	ram3 : Ram64
	port map(
		clock => clock,
		input => input,
		load => load,
		address => address( 5 downto 0),
		output => output
	);
	ram4 : Ram64
	port map(
		clock => clock,
		input => input,
		load => load,
		address => address( 5 downto 0),
		output => output
	);
	ram5 : Ram64
	port map(
		clock => clock,
		input => input,
		load => load,
		address => address( 5 downto 0),
		output => output
	);
	ram6 : Ram64
	port map(
		clock => clock,
		input => input,
		load => load,
		address => address( 5 downto 0),
		output => output
	);
	ram7 : Ram64
	port map(
		clock => clock,
		input => input,
		load => load,
		address => address( 5 downto 0),
		output => output
	);
end architecture;
