-- Elementos de Sistemas
-- FlipFlopJK.vhd

library ieee;
use ieee.std_logic_1164.all;

entity FlipFlopJK is
	port(
		clock:  in std_logic;
		J:      in std_logic;
		K:      in std_logic;
		q:      out std_logic:= '0';
		notq:   out std_logic:= '1'
	);
end entity;

architecture arch of FlipFlopJK is

signal q_conection, notq_conection : std_logic;

begin

	process (clock) begin
		if (rising_edge(clock) and J = '0' and K ='0') then
			q_conection <= q_conection;
			notq_conection <= notq_conection;
		elsif (rising_edge(clock) and J = '0' and K ='1') then
			q_conection <= '0';
			notq_conection <= '1';
		elsif (rising_edge(clock) and J = '1' and K ='0') then	
			q_conection <= '1';
			notq_conection <= '0';
		elsif (rising_edge(clock) and J = '1' and K ='1') then	
			q_conection <= notq_conection;
			notq_conection <= q_conection;
		end if;
	end process;
	q <= q_conection;
	notq <= notq_conection;
end architecture;
